//testbench for FFT_base2 module
`timescale 1ns / 1ps
module TB;





endmodule