//copyright (c) 2024 by LFQ
//email: lvfuq@outlook.com

//This module is used to generate the address for the FFT
